`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:44:22 10/21/2016 
// Design Name: 
// Module Name:    fft_128 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fft_128(
    input clk,
    input reset,
    input [15:0] re_in,
    input [15:0] im_in,
    output [15:0] re_out,
    output [15:0] im_out,
    input start,
    input valid_in,
    output valid_out
    );


endmodule
